//  -----------------------------------------------------------------------------
//                     Design Information
//  -----------------------------------------------------------------------------
//
//             Author: Begul Bilgin
//
//        Description: Mix Columns for the State
//
//  -----------------------------------------------------------------------------
module  mcol_state  ( a, y ) ;


input   [191:0]  a ;  // 4-bit input
output  [191:0]  y ;  // 4-bit yput

mcol m1(.a1(a[23:18]), .a2(a[17:12]), .a3(a[11:6]), .a4(a[5:0]), .y1(y[23:18]), .y2(y[17:12]), .y3(y[11:6]), .y4(y[5:0]) );
mcol m2(.a1(a[47:42]), .a2(a[41:36]), .a3(a[35:30]), .a4(a[29:24]), .y1(y[47:42]), .y2(y[41:36]), .y3(y[35:30]), .y4(y[29:24]) );
mcol m3(.a1(a[71:66]), .a2(a[65:60]), .a3(a[59:54]), .a4(a[53:48]), .y1(y[71:66]), .y2(y[65:60]), .y3(y[59:54]), .y4(y[53:48]) );
mcol m4(.a1(a[95:90]), .a2(a[89:84]), .a3(a[83:78]), .a4(a[77:72]), .y1(y[95:90]), .y2(y[89:84]), .y3(y[83:78]), .y4(y[77:72]) );
mcol m5(.a1(a[119:114]), .a2(a[113:108]), .a3(a[107:102]), .a4(a[101:96]), .y1(y[119:114]), .y2(y[113:108]), .y3(y[107:102]), .y4(y[101:96]) );
mcol m6(.a1(a[143:138]), .a2(a[137:132]), .a3(a[131:126]), .a4(a[125:120]), .y1(y[143:138]), .y2(y[137:132]), .y3(y[131:126]), .y4(y[125:120]) );
mcol m7(.a1(a[167:162]), .a2(a[161:156]), .a3(a[155:150]), .a4(a[149:144]), .y1(y[167:162]), .y2(y[161:156]), .y3(y[155:150]), .y4(y[149:144]) );
mcol m8(.a1(a[191:186]), .a2(a[185:180]), .a3(a[179:174]), .a4(a[173:168]), .y1(y[191:186]), .y2(y[185:180]), .y3(y[179:174]), .y4(y[173:168]) );


endmodule
