//  -----------------------------------------------------------------------------
//                     Design Information
//  -----------------------------------------------------------------------------
//
//             Author: Begul Bilgin
//
//        Description: 5-bit S-box, First Share File.
//
//  -----------------------------------------------------------------------------


//S:1   0  25  26  17  29  21  27  20   5   4  23  14  18   2  28  15   8   6   3  13   7  24  16  30   9  31  10  22  12  11  19

 module sbox_1 ( a2, a3, a4, y); 

input [0:4] a2; 
input [0:4] a3; 
input [0:4] a4; 
output [0:4] y; 

 assign y={a2[3]^a2[2]^((a2[3]^a3[3]^a4[3])&(a2[2]^a3[2]^a4[2]))^a2[1]^((a2[4]^a3[4]^a4[4])&(a2[1]^a3[1]^a4[1]))^((a2[3]^a3[3]^a4[3])&(a2[0]^a3[0]^a4[0]))^((a2[2]^a3[2]^a4[2])&(a2[0]^a3[0]^a4[0])),a2[3]^((a2[4]^a3[4]^a4[4])&(a2[2]^a3[2]^a4[2]))^((a2[3]^a3[3]^a4[3])&(a2[2]^a3[2]^a4[2]))^((a2[3]^a3[3]^a4[3])&(a2[1]^a3[1]^a4[1]))^((a2[2]^a3[2]^a4[2])&(a2[1]^a3[1]^a4[1]))^a2[0],((a2[4]^a3[4]^a4[4])&(a2[2]^a3[2]^a4[2]))^((a2[3]^a3[3]^a4[3])&(a2[2]^a3[2]^a4[2]))^a2[1]^a2[0]^((a2[4]^a3[4]^a4[4])&(a2[0]^a3[0]^a4[0]))^((a2[1]^a3[1]^a4[1])&(a2[0]^a3[0]^a4[0])),((a2[4]^a3[4]^a4[4])&(a2[3]^a3[3]^a4[3]))^((a2[2]^a3[2]^a4[2])&(a2[1]^a3[1]^a4[1]))^a2[0]^((a2[4]^a3[4]^a4[4])&(a2[0]^a3[0]^a4[0]))^((a2[2]^a3[2]^a4[2])&(a2[0]^a3[0]^a4[0])),1'b1^a2[4]^((a2[4]^a3[4]^a4[4])&(a2[2]^a3[2]^a4[2]))^a2[1]^((a2[3]^a3[3]^a4[3])&(a2[0]^a3[0]^a4[0]))}; 

 endmodule 
