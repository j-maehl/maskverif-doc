//  -----------------------------------------------------------------------------
//                     Design Information
//  -----------------------------------------------------------------------------
//
//             Author: Begul Bilgin
//
//        Description: 6-bit S-box for the State 
//
//  -----------------------------------------------------------------------------

 module sbox_state (a1,a2,a3,a4,y1,y2,y3,y4) ;

 input [191:0] a1;
 input [191:0] a2;
 input [191:0] a3;
 input [191:0] a4;
 output [191:0] y1;
 output [191:0] y2;
 output [191:0] y3;
 output [191:0] y4;
 
	f_1 sb01(.a2(a2[5:0]), .a3(a3[5:0]), .a4(a4[5:0]), .y(y1[5:0]));
	f_2 sb02(.a1(a1[5:0]), .a3(a3[5:0]), .a4(a4[5:0]), .y(y2[5:0]));
	f_3 sb03(.a1(a1[5:0]), .a2(a2[5:0]), .a4(a4[5:0]), .y(y3[5:0]));
	f_4 sb04(.a1(a1[5:0]), .a2(a2[5:0]), .a3(a3[5:0]), .y(y4[5:0]));

	f_1 sb11(.a2(a2[11:6]), .a3(a3[11:6]), .a4(a4[11:6]), .y(y1[11:6]));
	f_2 sb12(.a1(a1[11:6]), .a3(a3[11:6]), .a4(a4[11:6]), .y(y2[11:6]));
	f_3 sb13(.a1(a1[11:6]), .a2(a2[11:6]), .a4(a4[11:6]), .y(y3[11:6]));
	f_4 sb14(.a1(a1[11:6]), .a2(a2[11:6]), .a3(a3[11:6]), .y(y4[11:6]));

	f_1 sb21(.a2(a2[17:12]), .a3(a3[17:12]), .a4(a4[17:12]), .y(y1[17:12]));
	f_2 sb22(.a1(a1[17:12]), .a3(a3[17:12]), .a4(a4[17:12]), .y(y2[17:12]));
	f_3 sb23(.a1(a1[17:12]), .a2(a2[17:12]), .a4(a4[17:12]), .y(y3[17:12]));
	f_4 sb24(.a1(a1[17:12]), .a2(a2[17:12]), .a3(a3[17:12]), .y(y4[17:12]));

	f_1 sb31(.a2(a2[23:18]), .a3(a3[23:18]), .a4(a4[23:18]), .y(y1[23:18]));
	f_2 sb32(.a1(a1[23:18]), .a3(a3[23:18]), .a4(a4[23:18]), .y(y2[23:18]));
	f_3 sb33(.a1(a1[23:18]), .a2(a2[23:18]), .a4(a4[23:18]), .y(y3[23:18]));
	f_4 sb34(.a1(a1[23:18]), .a2(a2[23:18]), .a3(a3[23:18]), .y(y4[23:18]));

	f_1 sb41(.a2(a2[29:24]), .a3(a3[29:24]), .a4(a4[29:24]), .y(y1[29:24]));
	f_2 sb42(.a1(a1[29:24]), .a3(a3[29:24]), .a4(a4[29:24]), .y(y2[29:24]));
	f_3 sb43(.a1(a1[29:24]), .a2(a2[29:24]), .a4(a4[29:24]), .y(y3[29:24]));
	f_4 sb44(.a1(a1[29:24]), .a2(a2[29:24]), .a3(a3[29:24]), .y(y4[29:24]));

	f_1 sb51(.a2(a2[35:30]), .a3(a3[35:30]), .a4(a4[35:30]), .y(y1[35:30]));
	f_2 sb52(.a1(a1[35:30]), .a3(a3[35:30]), .a4(a4[35:30]), .y(y2[35:30]));
	f_3 sb53(.a1(a1[35:30]), .a2(a2[35:30]), .a4(a4[35:30]), .y(y3[35:30]));
	f_4 sb54(.a1(a1[35:30]), .a2(a2[35:30]), .a3(a3[35:30]), .y(y4[35:30]));

	f_1 sb61(.a2(a2[41:36]), .a3(a3[41:36]), .a4(a4[41:36]), .y(y1[41:36]));
	f_2 sb62(.a1(a1[41:36]), .a3(a3[41:36]), .a4(a4[41:36]), .y(y2[41:36]));
	f_3 sb63(.a1(a1[41:36]), .a2(a2[41:36]), .a4(a4[41:36]), .y(y3[41:36]));
	f_4 sb64(.a1(a1[41:36]), .a2(a2[41:36]), .a3(a3[41:36]), .y(y4[41:36]));

	f_1 sb71(.a2(a2[47:42]), .a3(a3[47:42]), .a4(a4[47:42]), .y(y1[47:42]));
	f_2 sb72(.a1(a1[47:42]), .a3(a3[47:42]), .a4(a4[47:42]), .y(y2[47:42]));
	f_3 sb73(.a1(a1[47:42]), .a2(a2[47:42]), .a4(a4[47:42]), .y(y3[47:42]));
	f_4 sb74(.a1(a1[47:42]), .a2(a2[47:42]), .a3(a3[47:42]), .y(y4[47:42]));

	f_1 sb81(.a2(a2[53:48]), .a3(a3[53:48]), .a4(a4[53:48]), .y(y1[53:48]));
	f_2 sb82(.a1(a1[53:48]), .a3(a3[53:48]), .a4(a4[53:48]), .y(y2[53:48]));
	f_3 sb83(.a1(a1[53:48]), .a2(a2[53:48]), .a4(a4[53:48]), .y(y3[53:48]));
	f_4 sb84(.a1(a1[53:48]), .a2(a2[53:48]), .a3(a3[53:48]), .y(y4[53:48]));

	f_1 sb91(.a2(a2[59:54]), .a3(a3[59:54]), .a4(a4[59:54]), .y(y1[59:54]));
	f_2 sb92(.a1(a1[59:54]), .a3(a3[59:54]), .a4(a4[59:54]), .y(y2[59:54]));
	f_3 sb93(.a1(a1[59:54]), .a2(a2[59:54]), .a4(a4[59:54]), .y(y3[59:54]));
	f_4 sb94(.a1(a1[59:54]), .a2(a2[59:54]), .a3(a3[59:54]), .y(y4[59:54]));

	f_1 sb101(.a2(a2[65:60]), .a3(a3[65:60]), .a4(a4[65:60]), .y(y1[65:60]));
	f_2 sb102(.a1(a1[65:60]), .a3(a3[65:60]), .a4(a4[65:60]), .y(y2[65:60]));
	f_3 sb103(.a1(a1[65:60]), .a2(a2[65:60]), .a4(a4[65:60]), .y(y3[65:60]));
	f_4 sb104(.a1(a1[65:60]), .a2(a2[65:60]), .a3(a3[65:60]), .y(y4[65:60]));

	f_1 sb111(.a2(a2[71:66]), .a3(a3[71:66]), .a4(a4[71:66]), .y(y1[71:66]));
	f_2 sb112(.a1(a1[71:66]), .a3(a3[71:66]), .a4(a4[71:66]), .y(y2[71:66]));
	f_3 sb113(.a1(a1[71:66]), .a2(a2[71:66]), .a4(a4[71:66]), .y(y3[71:66]));
	f_4 sb114(.a1(a1[71:66]), .a2(a2[71:66]), .a3(a3[71:66]), .y(y4[71:66]));

	f_1 sb121(.a2(a2[77:72]), .a3(a3[77:72]), .a4(a4[77:72]), .y(y1[77:72]));
	f_2 sb122(.a1(a1[77:72]), .a3(a3[77:72]), .a4(a4[77:72]), .y(y2[77:72]));
	f_3 sb123(.a1(a1[77:72]), .a2(a2[77:72]), .a4(a4[77:72]), .y(y3[77:72]));
	f_4 sb124(.a1(a1[77:72]), .a2(a2[77:72]), .a3(a3[77:72]), .y(y4[77:72]));

	f_1 sb131(.a2(a2[83:78]), .a3(a3[83:78]), .a4(a4[83:78]), .y(y1[83:78]));
	f_2 sb132(.a1(a1[83:78]), .a3(a3[83:78]), .a4(a4[83:78]), .y(y2[83:78]));
	f_3 sb133(.a1(a1[83:78]), .a2(a2[83:78]), .a4(a4[83:78]), .y(y3[83:78]));
	f_4 sb134(.a1(a1[83:78]), .a2(a2[83:78]), .a3(a3[83:78]), .y(y4[83:78]));

	f_1 sb141(.a2(a2[89:84]), .a3(a3[89:84]), .a4(a4[89:84]), .y(y1[89:84]));
	f_2 sb142(.a1(a1[89:84]), .a3(a3[89:84]), .a4(a4[89:84]), .y(y2[89:84]));
	f_3 sb143(.a1(a1[89:84]), .a2(a2[89:84]), .a4(a4[89:84]), .y(y3[89:84]));
	f_4 sb144(.a1(a1[89:84]), .a2(a2[89:84]), .a3(a3[89:84]), .y(y4[89:84]));

	f_1 sb151(.a2(a2[95:90]), .a3(a3[95:90]), .a4(a4[95:90]), .y(y1[95:90]));
	f_2 sb152(.a1(a1[95:90]), .a3(a3[95:90]), .a4(a4[95:90]), .y(y2[95:90]));
	f_3 sb153(.a1(a1[95:90]), .a2(a2[95:90]), .a4(a4[95:90]), .y(y3[95:90]));
	f_4 sb154(.a1(a1[95:90]), .a2(a2[95:90]), .a3(a3[95:90]), .y(y4[95:90]));

	f_1 sb161(.a2(a2[101:96]), .a3(a3[101:96]), .a4(a4[101:96]), .y(y1[101:96]));
	f_2 sb162(.a1(a1[101:96]), .a3(a3[101:96]), .a4(a4[101:96]), .y(y2[101:96]));
	f_3 sb163(.a1(a1[101:96]), .a2(a2[101:96]), .a4(a4[101:96]), .y(y3[101:96]));
	f_4 sb164(.a1(a1[101:96]), .a2(a2[101:96]), .a3(a3[101:96]), .y(y4[101:96]));

	f_1 sb171(.a2(a2[107:102]), .a3(a3[107:102]), .a4(a4[107:102]), .y(y1[107:102]));
	f_2 sb172(.a1(a1[107:102]), .a3(a3[107:102]), .a4(a4[107:102]), .y(y2[107:102]));
	f_3 sb173(.a1(a1[107:102]), .a2(a2[107:102]), .a4(a4[107:102]), .y(y3[107:102]));
	f_4 sb174(.a1(a1[107:102]), .a2(a2[107:102]), .a3(a3[107:102]), .y(y4[107:102]));

	f_1 sb181(.a2(a2[113:108]), .a3(a3[113:108]), .a4(a4[113:108]), .y(y1[113:108]));
	f_2 sb182(.a1(a1[113:108]), .a3(a3[113:108]), .a4(a4[113:108]), .y(y2[113:108]));
	f_3 sb183(.a1(a1[113:108]), .a2(a2[113:108]), .a4(a4[113:108]), .y(y3[113:108]));
	f_4 sb184(.a1(a1[113:108]), .a2(a2[113:108]), .a3(a3[113:108]), .y(y4[113:108]));

	f_1 sb191(.a2(a2[119:114]), .a3(a3[119:114]), .a4(a4[119:114]), .y(y1[119:114]));
	f_2 sb192(.a1(a1[119:114]), .a3(a3[119:114]), .a4(a4[119:114]), .y(y2[119:114]));
	f_3 sb193(.a1(a1[119:114]), .a2(a2[119:114]), .a4(a4[119:114]), .y(y3[119:114]));
	f_4 sb194(.a1(a1[119:114]), .a2(a2[119:114]), .a3(a3[119:114]), .y(y4[119:114]));

	f_1 sb201(.a2(a2[125:120]), .a3(a3[125:120]), .a4(a4[125:120]), .y(y1[125:120]));
	f_2 sb202(.a1(a1[125:120]), .a3(a3[125:120]), .a4(a4[125:120]), .y(y2[125:120]));
	f_3 sb203(.a1(a1[125:120]), .a2(a2[125:120]), .a4(a4[125:120]), .y(y3[125:120]));
	f_4 sb204(.a1(a1[125:120]), .a2(a2[125:120]), .a3(a3[125:120]), .y(y4[125:120]));

	f_1 sb211(.a2(a2[131:126]), .a3(a3[131:126]), .a4(a4[131:126]), .y(y1[131:126]));
	f_2 sb212(.a1(a1[131:126]), .a3(a3[131:126]), .a4(a4[131:126]), .y(y2[131:126]));
	f_3 sb213(.a1(a1[131:126]), .a2(a2[131:126]), .a4(a4[131:126]), .y(y3[131:126]));
	f_4 sb214(.a1(a1[131:126]), .a2(a2[131:126]), .a3(a3[131:126]), .y(y4[131:126]));

	f_1 sb221(.a2(a2[137:132]), .a3(a3[137:132]), .a4(a4[137:132]), .y(y1[137:132]));
	f_2 sb222(.a1(a1[137:132]), .a3(a3[137:132]), .a4(a4[137:132]), .y(y2[137:132]));
	f_3 sb223(.a1(a1[137:132]), .a2(a2[137:132]), .a4(a4[137:132]), .y(y3[137:132]));
	f_4 sb224(.a1(a1[137:132]), .a2(a2[137:132]), .a3(a3[137:132]), .y(y4[137:132]));

	f_1 sb231(.a2(a2[143:138]), .a3(a3[143:138]), .a4(a4[143:138]), .y(y1[143:138]));
	f_2 sb232(.a1(a1[143:138]), .a3(a3[143:138]), .a4(a4[143:138]), .y(y2[143:138]));
	f_3 sb233(.a1(a1[143:138]), .a2(a2[143:138]), .a4(a4[143:138]), .y(y3[143:138]));
	f_4 sb234(.a1(a1[143:138]), .a2(a2[143:138]), .a3(a3[143:138]), .y(y4[143:138]));

	f_1 sb241(.a2(a2[149:144]), .a3(a3[149:144]), .a4(a4[149:144]), .y(y1[149:144]));
	f_2 sb242(.a1(a1[149:144]), .a3(a3[149:144]), .a4(a4[149:144]), .y(y2[149:144]));
	f_3 sb243(.a1(a1[149:144]), .a2(a2[149:144]), .a4(a4[149:144]), .y(y3[149:144]));
	f_4 sb244(.a1(a1[149:144]), .a2(a2[149:144]), .a3(a3[149:144]), .y(y4[149:144]));

	f_1 sb251(.a2(a2[155:150]), .a3(a3[155:150]), .a4(a4[155:150]), .y(y1[155:150]));
	f_2 sb252(.a1(a1[155:150]), .a3(a3[155:150]), .a4(a4[155:150]), .y(y2[155:150]));
	f_3 sb253(.a1(a1[155:150]), .a2(a2[155:150]), .a4(a4[155:150]), .y(y3[155:150]));
	f_4 sb254(.a1(a1[155:150]), .a2(a2[155:150]), .a3(a3[155:150]), .y(y4[155:150]));

	f_1 sb261(.a2(a2[161:156]), .a3(a3[161:156]), .a4(a4[161:156]), .y(y1[161:156]));
	f_2 sb262(.a1(a1[161:156]), .a3(a3[161:156]), .a4(a4[161:156]), .y(y2[161:156]));
	f_3 sb263(.a1(a1[161:156]), .a2(a2[161:156]), .a4(a4[161:156]), .y(y3[161:156]));
	f_4 sb264(.a1(a1[161:156]), .a2(a2[161:156]), .a3(a3[161:156]), .y(y4[161:156]));

	f_1 sb271(.a2(a2[167:162]), .a3(a3[167:162]), .a4(a4[167:162]), .y(y1[167:162]));
	f_2 sb272(.a1(a1[167:162]), .a3(a3[167:162]), .a4(a4[167:162]), .y(y2[167:162]));
	f_3 sb273(.a1(a1[167:162]), .a2(a2[167:162]), .a4(a4[167:162]), .y(y3[167:162]));
	f_4 sb274(.a1(a1[167:162]), .a2(a2[167:162]), .a3(a3[167:162]), .y(y4[167:162]));

	f_1 sb281(.a2(a2[173:168]), .a3(a3[173:168]), .a4(a4[173:168]), .y(y1[173:168]));
	f_2 sb282(.a1(a1[173:168]), .a3(a3[173:168]), .a4(a4[173:168]), .y(y2[173:168]));
	f_3 sb283(.a1(a1[173:168]), .a2(a2[173:168]), .a4(a4[173:168]), .y(y3[173:168]));
	f_4 sb284(.a1(a1[173:168]), .a2(a2[173:168]), .a3(a3[173:168]), .y(y4[173:168]));

	f_1 sb291(.a2(a2[179:174]), .a3(a3[179:174]), .a4(a4[179:174]), .y(y1[179:174]));
	f_2 sb292(.a1(a1[179:174]), .a3(a3[179:174]), .a4(a4[179:174]), .y(y2[179:174]));
	f_3 sb293(.a1(a1[179:174]), .a2(a2[179:174]), .a4(a4[179:174]), .y(y3[179:174]));
	f_4 sb294(.a1(a1[179:174]), .a2(a2[179:174]), .a3(a3[179:174]), .y(y4[179:174]));

	f_1 sb301(.a2(a2[185:180]), .a3(a3[185:180]), .a4(a4[185:180]), .y(y1[185:180]));
	f_2 sb302(.a1(a1[185:180]), .a3(a3[185:180]), .a4(a4[185:180]), .y(y2[185:180]));
	f_3 sb303(.a1(a1[185:180]), .a2(a2[185:180]), .a4(a4[185:180]), .y(y3[185:180]));
	f_4 sb304(.a1(a1[185:180]), .a2(a2[185:180]), .a3(a3[185:180]), .y(y4[185:180]));

	f_1 sb311(.a2(a2[191:186]), .a3(a3[191:186]), .a4(a4[191:186]), .y(y1[191:186]));
	f_2 sb312(.a1(a1[191:186]), .a3(a3[191:186]), .a4(a4[191:186]), .y(y2[191:186]));
	f_3 sb313(.a1(a1[191:186]), .a2(a2[191:186]), .a4(a4[191:186]), .y(y3[191:186]));
	f_4 sb314(.a1(a1[191:186]), .a2(a2[191:186]), .a3(a3[191:186]), .y(y4[191:186]));
 endmodule 
