//  -----------------------------------------------------------------------------
//                     Design Information
//  -----------------------------------------------------------------------------
//
//             Author: Begul Bilgin
//
//        Description: Mix Columns for the State
//
//  -----------------------------------------------------------------------------
module  mcol_state  ( a, y ) ;


input   [159:0]  a ;  // 4-bit input

output  [159:0]  y ;  // 4-bit yput

wire [4:0] a00 = a[159:155];
wire [4:0] a01 = a[154:150];
wire [4:0] a02 = a[149:145];
wire [4:0] a03 = a[144:140];
wire [4:0] a10 = a[139:135];
wire [4:0] a11 = a[134:130];
wire [4:0] a12 = a[129:125];
wire [4:0] a13 = a[124:120];
wire [4:0] a20 = a[119:115];
wire [4:0] a21 = a[114:110];
wire [4:0] a22 = a[109:105];
wire [4:0] a23 = a[104:100];
wire [4:0] a30 = a[99:95];
wire [4:0] a31 = a[94:90];
wire [4:0] a32 = a[89:85];
wire [4:0] a33 = a[84:80];
wire [4:0] a40 = a[79:75];
wire [4:0] a41 = a[74:70];
wire [4:0] a42 = a[69:65];
wire [4:0] a43 = a[64:60];
wire [4:0] a50 = a[59:55];
wire [4:0] a51 = a[54:50];
wire [4:0] a52 = a[49:45];
wire [4:0] a53 = a[44:40];
wire [4:0] a60 = a[39:35];
wire [4:0] a61 = a[34:30];
wire [4:0] a62 = a[29:25];
wire [4:0] a63 = a[24:20];
wire [4:0] a70 = a[19:15];
wire [4:0] a71 = a[14:10];
wire [4:0] a72 = a[9:5];
wire [4:0] a73 = a[4:0];

mcol m1(.a1(a[159:155]), .a2(a[154:150]), .a3(a[149:145]), .a4(a[144:140]), .y1(y[159:155]), .y2(y[154:150]), .y3(y[149:145]), .y4(y[144:140]) );
mcol m2(.a1(a[139:135]), .a2(a[134:130]), .a3(a[129:125]), .a4(a[124:120]), .y1(y[139:135]), .y2(y[134:130]), .y3(y[129:125]), .y4(y[124:120]) );
mcol m3(.a1(a[119:115]), .a2(a[114:110]), .a3(a[109:105]), .a4(a[104:100]), .y1(y[119:115]), .y2(y[114:110]), .y3(y[109:105]), .y4(y[104:100]) );
mcol m4(.a1(a[99:95]), .a2(a[94:90]), .a3(a[89:85]), .a4(a[84:80]), .y1(y[99:95]), .y2(y[94:90]), .y3(y[89:85]), .y4(y[84:80]) );
mcol m5(.a1(a[79:75]), .a2(a[74:70]), .a3(a[69:65]), .a4(a[64:60]), .y1(y[79:75]), .y2(y[74:70]), .y3(y[69:65]), .y4(y[64:60]) );
mcol m6(.a1(a[59:55]), .a2(a[54:50]), .a3(a[49:45]), .a4(a[44:40]), .y1(y[59:55]), .y2(y[54:50]), .y3(y[49:45]), .y4(y[44:40]) );
mcol m7(.a1(a[39:35]), .a2(a[34:30]), .a3(a[29:25]), .a4(a[24:20]), .y1(y[39:35]), .y2(y[34:30]), .y3(y[29:25]), .y4(y[24:20]) );
mcol m8(.a1(a[19:15]), .a2(a[14:10]), .a3(a[9:5]), .a4(a[4:0]), .y1(y[19:15]), .y2(y[14:10]), .y3(y[9:5]), .y4(y[4:0]) );


endmodule
