//S:54   0  48  13  15  18  35  53  63  25  45  52   3  20  33  41   8  10  57  37  59  36  34   2  26  50  58  24  60  19  14  42  46  61   5  49  31  11  28   4  12  30  55  22   9   6  32  23  27  39  21  17  16  29  62   1  40  47  51  56   7  43  38  44

 module f_3 ( a1, a2, a4, y); 

input [0:5] a1; 
input [0:5] a2; 
input [0:5] a4; 
output [0:5] y; 

 assign y={a4[5]^a4[3]^(a1[5]&a2[3])^(a2[5]&a1[3])^(a1[4]&a2[3])^(a2[4]&a1[3])^(a1[2]&a1[4]&a2[5])^(a1[2]&a2[4]&a1[5])^(a2[2]&a1[4]&a1[5])^(a1[2]&a2[4]&a2[5])^(a2[2]&a1[4]&a2[5])^(a2[2]&a2[4]&a1[5])^(a1[2]&a2[4]&a4[5])^(a2[2]&a1[4]&a4[5])^(a1[2]&a4[4]&a2[5])^(a2[2]&a4[4]&a1[5])^(a4[2]&a1[4]&a2[5])^(a4[2]&a2[4]&a1[5])^a4[1]^(a1[5]&a2[1])^(a2[5]&a1[1])^(a1[4]&a2[1])^(a2[4]&a1[1])^(a1[1]&a1[3]&a2[5])^(a1[1]&a2[3]&a1[5])^(a2[1]&a1[3]&a1[5])^(a1[1]&a2[3]&a2[5])^(a2[1]&a1[3]&a2[5])^(a2[1]&a2[3]&a1[5])^(a1[1]&a2[3]&a4[5])^(a2[1]&a1[3]&a4[5])^(a1[1]&a4[3]&a2[5])^(a2[1]&a4[3]&a1[5])^(a4[1]&a1[3]&a2[5])^(a4[1]&a2[3]&a1[5])^(a1[1]&a1[2]&a2[5])^(a1[1]&a2[2]&a1[5])^(a2[1]&a1[2]&a1[5])^(a1[1]&a2[2]&a2[5])^(a2[1]&a1[2]&a2[5])^(a2[1]&a2[2]&a1[5])^(a1[1]&a2[2]&a4[5])^(a2[1]&a1[2]&a4[5])^(a1[1]&a4[2]&a2[5])^(a2[1]&a4[2]&a1[5])^(a4[1]&a1[2]&a2[5])^(a4[1]&a2[2]&a1[5])^(a1[5]&a2[0])^(a2[5]&a1[0])^(a1[4]&a2[0])^(a2[4]&a1[0])^(a1[0]&a1[4]&a2[5])^(a1[0]&a2[4]&a1[5])^(a2[0]&a1[4]&a1[5])^(a1[0]&a2[4]&a2[5])^(a2[0]&a1[4]&a2[5])^(a2[0]&a2[4]&a1[5])^(a1[0]&a2[4]&a4[5])^(a2[0]&a1[4]&a4[5])^(a1[0]&a4[4]&a2[5])^(a2[0]&a4[4]&a1[5])^(a4[0]&a1[4]&a2[5])^(a4[0]&a2[4]&a1[5])^(a1[0]&a1[3]&a2[5])^(a1[0]&a2[3]&a1[5])^(a2[0]&a1[3]&a1[5])^(a1[0]&a2[3]&a2[5])^(a2[0]&a1[3]&a2[5])^(a2[0]&a2[3]&a1[5])^(a1[0]&a2[3]&a4[5])^(a2[0]&a1[3]&a4[5])^(a1[0]&a4[3]&a2[5])^(a2[0]&a4[3]&a1[5])^(a4[0]&a1[3]&a2[5])^(a4[0]&a2[3]&a1[5])^(a1[2]&a2[0])^(a2[2]&a1[0])^(a1[0]&a1[2]&a2[3])^(a1[0]&a2[2]&a1[3])^(a2[0]&a1[2]&a1[3])^(a1[0]&a2[2]&a2[3])^(a2[0]&a1[2]&a2[3])^(a2[0]&a2[2]&a1[3])^(a1[0]&a2[2]&a4[3])^(a2[0]&a1[2]&a4[3])^(a1[0]&a4[2]&a2[3])^(a2[0]&a4[2]&a1[3])^(a4[0]&a1[2]&a2[3])^(a4[0]&a2[2]&a1[3])^(a1[0]&a1[1]&a2[3])^(a1[0]&a2[1]&a1[3])^(a2[0]&a1[1]&a1[3])^(a1[0]&a2[1]&a2[3])^(a2[0]&a1[1]&a2[3])^(a2[0]&a2[1]&a1[3])^(a1[0]&a2[1]&a4[3])^(a2[0]&a1[1]&a4[3])^(a1[0]&a4[1]&a2[3])^(a2[0]&a4[1]&a1[3])^(a4[0]&a1[1]&a2[3])^(a4[0]&a2[1]&a1[3]),a4[5]^a4[3]^(a1[5]&a2[2])^(a2[5]&a1[2])^(a1[4]&a2[2])^(a2[4]&a1[2])^(a1[2]&a1[4]&a2[5])^(a1[2]&a2[4]&a1[5])^(a2[2]&a1[4]&a1[5])^(a1[2]&a2[4]&a2[5])^(a2[2]&a1[4]&a2[5])^(a2[2]&a2[4]&a1[5])^(a1[2]&a2[4]&a4[5])^(a2[2]&a1[4]&a4[5])^(a1[2]&a4[4]&a2[5])^(a2[2]&a4[4]&a1[5])^(a4[2]&a1[4]&a2[5])^(a4[2]&a2[4]&a1[5])^(a1[2]&a1[3]&a2[5])^(a1[2]&a2[3]&a1[5])^(a2[2]&a1[3]&a1[5])^(a1[2]&a2[3]&a2[5])^(a2[2]&a1[3]&a2[5])^(a2[2]&a2[3]&a1[5])^(a1[2]&a2[3]&a4[5])^(a2[2]&a1[3]&a4[5])^(a1[2]&a4[3]&a2[5])^(a2[2]&a4[3]&a1[5])^(a4[2]&a1[3]&a2[5])^(a4[2]&a2[3]&a1[5])^(a1[2]&a1[3]&a2[4])^(a1[2]&a2[3]&a1[4])^(a2[2]&a1[3]&a1[4])^(a1[2]&a2[3]&a2[4])^(a2[2]&a1[3]&a2[4])^(a2[2]&a2[3]&a1[4])^(a1[2]&a2[3]&a4[4])^(a2[2]&a1[3]&a4[4])^(a1[2]&a4[3]&a2[4])^(a2[2]&a4[3]&a1[4])^(a4[2]&a1[3]&a2[4])^(a4[2]&a2[3]&a1[4])^a4[1]^(a1[5]&a2[1])^(a2[5]&a1[1])^(a1[4]&a2[1])^(a2[4]&a1[1])^(a1[1]&a1[4]&a2[5])^(a1[1]&a2[4]&a1[5])^(a2[1]&a1[4]&a1[5])^(a1[1]&a2[4]&a2[5])^(a2[1]&a1[4]&a2[5])^(a2[1]&a2[4]&a1[5])^(a1[1]&a2[4]&a4[5])^(a2[1]&a1[4]&a4[5])^(a1[1]&a4[4]&a2[5])^(a2[1]&a4[4]&a1[5])^(a4[1]&a1[4]&a2[5])^(a4[1]&a2[4]&a1[5])^(a1[1]&a1[3]&a2[5])^(a1[1]&a2[3]&a1[5])^(a2[1]&a1[3]&a1[5])^(a1[1]&a2[3]&a2[5])^(a2[1]&a1[3]&a2[5])^(a2[1]&a2[3]&a1[5])^(a1[1]&a2[3]&a4[5])^(a2[1]&a1[3]&a4[5])^(a1[1]&a4[3]&a2[5])^(a2[1]&a4[3]&a1[5])^(a4[1]&a1[3]&a2[5])^(a4[1]&a2[3]&a1[5])^(a1[2]&a2[1])^(a2[2]&a1[1])^(a1[1]&a1[2]&a2[5])^(a1[1]&a2[2]&a1[5])^(a2[1]&a1[2]&a1[5])^(a1[1]&a2[2]&a2[5])^(a2[1]&a1[2]&a2[5])^(a2[1]&a2[2]&a1[5])^(a1[1]&a2[2]&a4[5])^(a2[1]&a1[2]&a4[5])^(a1[1]&a4[2]&a2[5])^(a2[1]&a4[2]&a1[5])^(a4[1]&a1[2]&a2[5])^(a4[1]&a2[2]&a1[5])^(a1[1]&a1[2]&a2[3])^(a1[1]&a2[2]&a1[3])^(a2[1]&a1[2]&a1[3])^(a1[1]&a2[2]&a2[3])^(a2[1]&a1[2]&a2[3])^(a2[1]&a2[2]&a1[3])^(a1[1]&a2[2]&a4[3])^(a2[1]&a1[2]&a4[3])^(a1[1]&a4[2]&a2[3])^(a2[1]&a4[2]&a1[3])^(a4[1]&a1[2]&a2[3])^(a4[1]&a2[2]&a1[3])^a4[0]^(a1[0]&a1[2]&a2[5])^(a1[0]&a2[2]&a1[5])^(a2[0]&a1[2]&a1[5])^(a1[0]&a2[2]&a2[5])^(a2[0]&a1[2]&a2[5])^(a2[0]&a2[2]&a1[5])^(a1[0]&a2[2]&a4[5])^(a2[0]&a1[2]&a4[5])^(a1[0]&a4[2]&a2[5])^(a2[0]&a4[2]&a1[5])^(a4[0]&a1[2]&a2[5])^(a4[0]&a2[2]&a1[5])^(a1[0]&a1[2]&a2[3])^(a1[0]&a2[2]&a1[3])^(a2[0]&a1[2]&a1[3])^(a1[0]&a2[2]&a2[3])^(a2[0]&a1[2]&a2[3])^(a2[0]&a2[2]&a1[3])^(a1[0]&a2[2]&a4[3])^(a2[0]&a1[2]&a4[3])^(a1[0]&a4[2]&a2[3])^(a2[0]&a4[2]&a1[3])^(a4[0]&a1[2]&a2[3])^(a4[0]&a2[2]&a1[3])^(a1[0]&a1[1]&a2[5])^(a1[0]&a2[1]&a1[5])^(a2[0]&a1[1]&a1[5])^(a1[0]&a2[1]&a2[5])^(a2[0]&a1[1]&a2[5])^(a2[0]&a2[1]&a1[5])^(a1[0]&a2[1]&a4[5])^(a2[0]&a1[1]&a4[5])^(a1[0]&a4[1]&a2[5])^(a2[0]&a4[1]&a1[5])^(a4[0]&a1[1]&a2[5])^(a4[0]&a2[1]&a1[5])^(a1[0]&a1[1]&a2[4])^(a1[0]&a2[1]&a1[4])^(a2[0]&a1[1]&a1[4])^(a1[0]&a2[1]&a2[4])^(a2[0]&a1[1]&a2[4])^(a2[0]&a2[1]&a1[4])^(a1[0]&a2[1]&a4[4])^(a2[0]&a1[1]&a4[4])^(a1[0]&a4[1]&a2[4])^(a2[0]&a4[1]&a1[4])^(a4[0]&a1[1]&a2[4])^(a4[0]&a2[1]&a1[4])^(a1[0]&a1[1]&a2[3])^(a1[0]&a2[1]&a1[3])^(a2[0]&a1[1]&a1[3])^(a1[0]&a2[1]&a2[3])^(a2[0]&a1[1]&a2[3])^(a2[0]&a2[1]&a1[3])^(a1[0]&a2[1]&a4[3])^(a2[0]&a1[1]&a4[3])^(a1[0]&a4[1]&a2[3])^(a2[0]&a4[1]&a1[3])^(a4[0]&a1[1]&a2[3])^(a4[0]&a2[1]&a1[3]),(a1[5]&a2[4])^(a2[5]&a1[4])^a4[3]^(a1[5]&a2[3])^(a2[5]&a1[3])^(a1[4]&a2[3])^(a2[4]&a1[3])^a4[2]^(a1[2]&a1[3]&a2[5])^(a1[2]&a2[3]&a1[5])^(a2[2]&a1[3]&a1[5])^(a1[2]&a2[3]&a2[5])^(a2[2]&a1[3]&a2[5])^(a2[2]&a2[3]&a1[5])^(a1[2]&a2[3]&a4[5])^(a2[2]&a1[3]&a4[5])^(a1[2]&a4[3]&a2[5])^(a2[2]&a4[3]&a1[5])^(a4[2]&a1[3]&a2[5])^(a4[2]&a2[3]&a1[5])^(a1[2]&a1[3]&a2[4])^(a1[2]&a2[3]&a1[4])^(a2[2]&a1[3]&a1[4])^(a1[2]&a2[3]&a2[4])^(a2[2]&a1[3]&a2[4])^(a2[2]&a2[3]&a1[4])^(a1[2]&a2[3]&a4[4])^(a2[2]&a1[3]&a4[4])^(a1[2]&a4[3]&a2[4])^(a2[2]&a4[3]&a1[4])^(a4[2]&a1[3]&a2[4])^(a4[2]&a2[3]&a1[4])^a4[1]^(a1[3]&a2[1])^(a2[3]&a1[1])^(a1[2]&a2[1])^(a2[2]&a1[1])^(a1[1]&a1[2]&a2[5])^(a1[1]&a2[2]&a1[5])^(a2[1]&a1[2]&a1[5])^(a1[1]&a2[2]&a2[5])^(a2[1]&a1[2]&a2[5])^(a2[1]&a2[2]&a1[5])^(a1[1]&a2[2]&a4[5])^(a2[1]&a1[2]&a4[5])^(a1[1]&a4[2]&a2[5])^(a2[1]&a4[2]&a1[5])^(a4[1]&a1[2]&a2[5])^(a4[1]&a2[2]&a1[5])^a4[0]^(a1[4]&a2[0])^(a2[4]&a1[0])^(a1[0]&a1[4]&a2[5])^(a1[0]&a2[4]&a1[5])^(a2[0]&a1[4]&a1[5])^(a1[0]&a2[4]&a2[5])^(a2[0]&a1[4]&a2[5])^(a2[0]&a2[4]&a1[5])^(a1[0]&a2[4]&a4[5])^(a2[0]&a1[4]&a4[5])^(a1[0]&a4[4]&a2[5])^(a2[0]&a4[4]&a1[5])^(a4[0]&a1[4]&a2[5])^(a4[0]&a2[4]&a1[5])^(a1[3]&a2[0])^(a2[3]&a1[0])^(a1[0]&a1[3]&a2[5])^(a1[0]&a2[3]&a1[5])^(a2[0]&a1[3]&a1[5])^(a1[0]&a2[3]&a2[5])^(a2[0]&a1[3]&a2[5])^(a2[0]&a2[3]&a1[5])^(a1[0]&a2[3]&a4[5])^(a2[0]&a1[3]&a4[5])^(a1[0]&a4[3]&a2[5])^(a2[0]&a4[3]&a1[5])^(a4[0]&a1[3]&a2[5])^(a4[0]&a2[3]&a1[5])^(a1[2]&a2[0])^(a2[2]&a1[0])^(a1[1]&a2[0])^(a2[1]&a1[0])^(a1[0]&a1[1]&a2[5])^(a1[0]&a2[1]&a1[5])^(a2[0]&a1[1]&a1[5])^(a1[0]&a2[1]&a2[5])^(a2[0]&a1[1]&a2[5])^(a2[0]&a2[1]&a1[5])^(a1[0]&a2[1]&a4[5])^(a2[0]&a1[1]&a4[5])^(a1[0]&a4[1]&a2[5])^(a2[0]&a4[1]&a1[5])^(a4[0]&a1[1]&a2[5])^(a4[0]&a2[1]&a1[5])^(a1[0]&a1[1]&a2[2])^(a1[0]&a2[1]&a1[2])^(a2[0]&a1[1]&a1[2])^(a1[0]&a2[1]&a2[2])^(a2[0]&a1[1]&a2[2])^(a2[0]&a2[1]&a1[2])^(a1[0]&a2[1]&a4[2])^(a2[0]&a1[1]&a4[2])^(a1[0]&a4[1]&a2[2])^(a2[0]&a4[1]&a1[2])^(a4[0]&a1[1]&a2[2])^(a4[0]&a2[1]&a1[2]),a4[5]^a4[4]^(a1[4]&a2[2])^(a2[4]&a1[2])^(a1[2]&a1[4]&a2[5])^(a1[2]&a2[4]&a1[5])^(a2[2]&a1[4]&a1[5])^(a1[2]&a2[4]&a2[5])^(a2[2]&a1[4]&a2[5])^(a2[2]&a2[4]&a1[5])^(a1[2]&a2[4]&a4[5])^(a2[2]&a1[4]&a4[5])^(a1[2]&a4[4]&a2[5])^(a2[2]&a4[4]&a1[5])^(a4[2]&a1[4]&a2[5])^(a4[2]&a2[4]&a1[5])^(a1[3]&a2[2])^(a2[3]&a1[2])^a4[1]^(a1[5]&a2[1])^(a2[5]&a1[1])^(a1[4]&a2[1])^(a2[4]&a1[1])^(a1[1]&a1[4]&a2[5])^(a1[1]&a2[4]&a1[5])^(a2[1]&a1[4]&a1[5])^(a1[1]&a2[4]&a2[5])^(a2[1]&a1[4]&a2[5])^(a2[1]&a2[4]&a1[5])^(a1[1]&a2[4]&a4[5])^(a2[1]&a1[4]&a4[5])^(a1[1]&a4[4]&a2[5])^(a2[1]&a4[4]&a1[5])^(a4[1]&a1[4]&a2[5])^(a4[1]&a2[4]&a1[5])^(a1[1]&a1[3]&a2[5])^(a1[1]&a2[3]&a1[5])^(a2[1]&a1[3]&a1[5])^(a1[1]&a2[3]&a2[5])^(a2[1]&a1[3]&a2[5])^(a2[1]&a2[3]&a1[5])^(a1[1]&a2[3]&a4[5])^(a2[1]&a1[3]&a4[5])^(a1[1]&a4[3]&a2[5])^(a2[1]&a4[3]&a1[5])^(a4[1]&a1[3]&a2[5])^(a4[1]&a2[3]&a1[5])^(a1[1]&a1[2]&a2[4])^(a1[1]&a2[2]&a1[4])^(a2[1]&a1[2]&a1[4])^(a1[1]&a2[2]&a2[4])^(a2[1]&a1[2]&a2[4])^(a2[1]&a2[2]&a1[4])^(a1[1]&a2[2]&a4[4])^(a2[1]&a1[2]&a4[4])^(a1[1]&a4[2]&a2[4])^(a2[1]&a4[2]&a1[4])^(a4[1]&a1[2]&a2[4])^(a4[1]&a2[2]&a1[4])^(a1[5]&a2[0])^(a2[5]&a1[0])^(a1[4]&a2[0])^(a2[4]&a1[0])^(a1[0]&a1[4]&a2[5])^(a1[0]&a2[4]&a1[5])^(a2[0]&a1[4]&a1[5])^(a1[0]&a2[4]&a2[5])^(a2[0]&a1[4]&a2[5])^(a2[0]&a2[4]&a1[5])^(a1[0]&a2[4]&a4[5])^(a2[0]&a1[4]&a4[5])^(a1[0]&a4[4]&a2[5])^(a2[0]&a4[4]&a1[5])^(a4[0]&a1[4]&a2[5])^(a4[0]&a2[4]&a1[5])^(a1[0]&a1[3]&a2[5])^(a1[0]&a2[3]&a1[5])^(a2[0]&a1[3]&a1[5])^(a1[0]&a2[3]&a2[5])^(a2[0]&a1[3]&a2[5])^(a2[0]&a2[3]&a1[5])^(a1[0]&a2[3]&a4[5])^(a2[0]&a1[3]&a4[5])^(a1[0]&a4[3]&a2[5])^(a2[0]&a4[3]&a1[5])^(a4[0]&a1[3]&a2[5])^(a4[0]&a2[3]&a1[5])^(a1[0]&a1[2]&a2[4])^(a1[0]&a2[2]&a1[4])^(a2[0]&a1[2]&a1[4])^(a1[0]&a2[2]&a2[4])^(a2[0]&a1[2]&a2[4])^(a2[0]&a2[2]&a1[4])^(a1[0]&a2[2]&a4[4])^(a2[0]&a1[2]&a4[4])^(a1[0]&a4[2]&a2[4])^(a2[0]&a4[2]&a1[4])^(a4[0]&a1[2]&a2[4])^(a4[0]&a2[2]&a1[4]),a4[5]^a4[4]^(a1[5]&a2[4])^(a2[5]&a1[4])^(a1[5]&a2[3])^(a2[5]&a1[3])^(a1[4]&a2[3])^(a2[4]&a1[3])^(a1[2]&a1[3]&a2[5])^(a1[2]&a2[3]&a1[5])^(a2[2]&a1[3]&a1[5])^(a1[2]&a2[3]&a2[5])^(a2[2]&a1[3]&a2[5])^(a2[2]&a2[3]&a1[5])^(a1[2]&a2[3]&a4[5])^(a2[2]&a1[3]&a4[5])^(a1[2]&a4[3]&a2[5])^(a2[2]&a4[3]&a1[5])^(a4[2]&a1[3]&a2[5])^(a4[2]&a2[3]&a1[5])^(a1[2]&a1[3]&a2[4])^(a1[2]&a2[3]&a1[4])^(a2[2]&a1[3]&a1[4])^(a1[2]&a2[3]&a2[4])^(a2[2]&a1[3]&a2[4])^(a2[2]&a2[3]&a1[4])^(a1[2]&a2[3]&a4[4])^(a2[2]&a1[3]&a4[4])^(a1[2]&a4[3]&a2[4])^(a2[2]&a4[3]&a1[4])^(a4[2]&a1[3]&a2[4])^(a4[2]&a2[3]&a1[4])^a4[1]^(a1[4]&a2[1])^(a2[4]&a1[1])^(a1[3]&a2[1])^(a2[3]&a1[1])^(a1[1]&a1[3]&a2[5])^(a1[1]&a2[3]&a1[5])^(a2[1]&a1[3]&a1[5])^(a1[1]&a2[3]&a2[5])^(a2[1]&a1[3]&a2[5])^(a2[1]&a2[3]&a1[5])^(a1[1]&a2[3]&a4[5])^(a2[1]&a1[3]&a4[5])^(a1[1]&a4[3]&a2[5])^(a2[1]&a4[3]&a1[5])^(a4[1]&a1[3]&a2[5])^(a4[1]&a2[3]&a1[5])^(a1[1]&a1[3]&a2[4])^(a1[1]&a2[3]&a1[4])^(a2[1]&a1[3]&a1[4])^(a1[1]&a2[3]&a2[4])^(a2[1]&a1[3]&a2[4])^(a2[1]&a2[3]&a1[4])^(a1[1]&a2[3]&a4[4])^(a2[1]&a1[3]&a4[4])^(a1[1]&a4[3]&a2[4])^(a2[1]&a4[3]&a1[4])^(a4[1]&a1[3]&a2[4])^(a4[1]&a2[3]&a1[4])^(a1[2]&a2[1])^(a2[2]&a1[1])^(a1[1]&a1[2]&a2[5])^(a1[1]&a2[2]&a1[5])^(a2[1]&a1[2]&a1[5])^(a1[1]&a2[2]&a2[5])^(a2[1]&a1[2]&a2[5])^(a2[1]&a2[2]&a1[5])^(a1[1]&a2[2]&a4[5])^(a2[1]&a1[2]&a4[5])^(a1[1]&a4[2]&a2[5])^(a2[1]&a4[2]&a1[5])^(a4[1]&a1[2]&a2[5])^(a4[1]&a2[2]&a1[5])^(a1[0]&a1[3]&a2[4])^(a1[0]&a2[3]&a1[4])^(a2[0]&a1[3]&a1[4])^(a1[0]&a2[3]&a2[4])^(a2[0]&a1[3]&a2[4])^(a2[0]&a2[3]&a1[4])^(a1[0]&a2[3]&a4[4])^(a2[0]&a1[3]&a4[4])^(a1[0]&a4[3]&a2[4])^(a2[0]&a4[3]&a1[4])^(a4[0]&a1[3]&a2[4])^(a4[0]&a2[3]&a1[4])^(a1[2]&a2[0])^(a2[2]&a1[0])^(a1[1]&a2[0])^(a2[1]&a1[0])^(a1[0]&a1[1]&a2[5])^(a1[0]&a2[1]&a1[5])^(a2[0]&a1[1]&a1[5])^(a1[0]&a2[1]&a2[5])^(a2[0]&a1[1]&a2[5])^(a2[0]&a2[1]&a1[5])^(a1[0]&a2[1]&a4[5])^(a2[0]&a1[1]&a4[5])^(a1[0]&a4[1]&a2[5])^(a2[0]&a4[1]&a1[5])^(a4[0]&a1[1]&a2[5])^(a4[0]&a2[1]&a1[5])^(a1[0]&a1[1]&a2[4])^(a1[0]&a2[1]&a1[4])^(a2[0]&a1[1]&a1[4])^(a1[0]&a2[1]&a2[4])^(a2[0]&a1[1]&a2[4])^(a2[0]&a2[1]&a1[4])^(a1[0]&a2[1]&a4[4])^(a2[0]&a1[1]&a4[4])^(a1[0]&a4[1]&a2[4])^(a2[0]&a4[1]&a1[4])^(a4[0]&a1[1]&a2[4])^(a4[0]&a2[1]&a1[4])^(a1[0]&a1[1]&a2[2])^(a1[0]&a2[1]&a1[2])^(a2[0]&a1[1]&a1[2])^(a1[0]&a2[1]&a2[2])^(a2[0]&a1[1]&a2[2])^(a2[0]&a2[1]&a1[2])^(a1[0]&a2[1]&a4[2])^(a2[0]&a1[1]&a4[2])^(a1[0]&a4[1]&a2[2])^(a2[0]&a4[1]&a1[2])^(a4[0]&a1[1]&a2[2])^(a4[0]&a2[1]&a1[2]),(a1[5]&a2[4])^(a2[5]&a1[4])^a4[3]^(a1[5]&a2[3])^(a2[5]&a1[3])^a4[2]^(a1[3]&a2[2])^(a2[3]&a1[2])^(a1[4]&a2[1])^(a2[4]&a1[1])^(a1[1]&a1[4]&a2[5])^(a1[1]&a2[4]&a1[5])^(a2[1]&a1[4]&a1[5])^(a1[1]&a2[4]&a2[5])^(a2[1]&a1[4]&a2[5])^(a2[1]&a2[4]&a1[5])^(a1[1]&a2[4]&a4[5])^(a2[1]&a1[4]&a4[5])^(a1[1]&a4[4]&a2[5])^(a2[1]&a4[4]&a1[5])^(a4[1]&a1[4]&a2[5])^(a4[1]&a2[4]&a1[5])^(a1[2]&a2[1])^(a2[2]&a1[1])^(a1[1]&a1[2]&a2[4])^(a1[1]&a2[2]&a1[4])^(a2[1]&a1[2]&a1[4])^(a1[1]&a2[2]&a2[4])^(a2[1]&a1[2]&a2[4])^(a2[1]&a2[2]&a1[4])^(a1[1]&a2[2]&a4[4])^(a2[1]&a1[2]&a4[4])^(a1[1]&a4[2]&a2[4])^(a2[1]&a4[2]&a1[4])^(a4[1]&a1[2]&a2[4])^(a4[1]&a2[2]&a1[4])^(a1[5]&a2[0])^(a2[5]&a1[0])^(a1[4]&a2[0])^(a2[4]&a1[0])^(a1[2]&a2[0])^(a2[2]&a1[0])^(a1[0]&a1[2]&a2[5])^(a1[0]&a2[2]&a1[5])^(a2[0]&a1[2]&a1[5])^(a1[0]&a2[2]&a2[5])^(a2[0]&a1[2]&a2[5])^(a2[0]&a2[2]&a1[5])^(a1[0]&a2[2]&a4[5])^(a2[0]&a1[2]&a4[5])^(a1[0]&a4[2]&a2[5])^(a2[0]&a4[2]&a1[5])^(a4[0]&a1[2]&a2[5])^(a4[0]&a2[2]&a1[5])^(a1[0]&a1[2]&a2[3])^(a1[0]&a2[2]&a1[3])^(a2[0]&a1[2]&a1[3])^(a1[0]&a2[2]&a2[3])^(a2[0]&a1[2]&a2[3])^(a2[0]&a2[2]&a1[3])^(a1[0]&a2[2]&a4[3])^(a2[0]&a1[2]&a4[3])^(a1[0]&a4[2]&a2[3])^(a2[0]&a4[2]&a1[3])^(a4[0]&a1[2]&a2[3])^(a4[0]&a2[2]&a1[3])^(a1[1]&a2[0])^(a2[1]&a1[0])^(a1[0]&a1[1]&a2[5])^(a1[0]&a2[1]&a1[5])^(a2[0]&a1[1]&a1[5])^(a1[0]&a2[1]&a2[5])^(a2[0]&a1[1]&a2[5])^(a2[0]&a2[1]&a1[5])^(a1[0]&a2[1]&a4[5])^(a2[0]&a1[1]&a4[5])^(a1[0]&a4[1]&a2[5])^(a2[0]&a4[1]&a1[5])^(a4[0]&a1[1]&a2[5])^(a4[0]&a2[1]&a1[5])}; 

 endmodule 
