//  -----------------------------------------------------------------------------
//                     Design Information
//  -----------------------------------------------------------------------------
//
//             Author: Begul Bilgin
//
//        Description: 5-bit S-box, Fourth Share File.
//
//  -----------------------------------------------------------------------------

//S:1   0  25  26  17  29  21  27  20   5   4  23  14  18   2  28  15   8   6   3  13   7  24  16  30   9  31  10  22  12  11  19

 module sbox_4 ( a1, a2, a3, y); 

input [0:4] a1; 
input [0:4] a2; 
input [0:4] a3; 
output [0:4] y; 

 assign y={a1[3]^a1[2]^a1[1],a1[3]^a1[0],a1[1]^a1[0],a1[0],a1[4]^a1[1]}; 

 endmodule 
