//  -----------------------------------------------------------------------------
//                     Design Information
//  -----------------------------------------------------------------------------
//
//             Author: Begul Bilgin
//
//        Description: 5-bit S-box for the State 
//
//  -----------------------------------------------------------------------------

//5x5 Sbox 
//S:1   0  25  26  17  29  21  27  20   5   4  23  14  18   2  28  15   8   6   3  13   7  24  16  30   9  31  10  22  12  11  19

 module sbox_state (a1,a2,a3,a4,y1,y2,y3,y4) ;

 input [159:0] a1;
 input [159:0] a2;
 input [159:0] a3;
 input [159:0] a4;
 output [159:0] y1;
 output [159:0] y2;
 output [159:0] y3;
 output [159:0] y4;
 
	sbox_1 sb01(.a2(a2[4:0]), .a3(a3[4:0]), .a4(a4[4:0]), .y(y1[4:0]));
	sbox_2 sb02(.a1(a1[4:0]), .a3(a3[4:0]), .a4(a4[4:0]), .y(y2[4:0]));
	sbox_3 sb03(.a1(a1[4:0]), .a2(a2[4:0]), .a4(a4[4:0]), .y(y3[4:0]));
	sbox_4 sb04(.a1(a1[4:0]), .a2(a2[4:0]), .a3(a3[4:0]), .y(y4[4:0]));

	sbox_1 sb11(.a2(a2[9:5]), .a3(a3[9:5]), .a4(a4[9:5]), .y(y1[9:5]));
	sbox_2 sb12(.a1(a1[9:5]), .a3(a3[9:5]), .a4(a4[9:5]), .y(y2[9:5]));
	sbox_3 sb13(.a1(a1[9:5]), .a2(a2[9:5]), .a4(a4[9:5]), .y(y3[9:5]));
	sbox_4 sb14(.a1(a1[9:5]), .a2(a2[9:5]), .a3(a3[9:5]), .y(y4[9:5]));

	sbox_1 sb21(.a2(a2[14:10]), .a3(a3[14:10]), .a4(a4[14:10]), .y(y1[14:10]));
	sbox_2 sb22(.a1(a1[14:10]), .a3(a3[14:10]), .a4(a4[14:10]), .y(y2[14:10]));
	sbox_3 sb23(.a1(a1[14:10]), .a2(a2[14:10]), .a4(a4[14:10]), .y(y3[14:10]));
	sbox_4 sb24(.a1(a1[14:10]), .a2(a2[14:10]), .a3(a3[14:10]), .y(y4[14:10]));

	sbox_1 sb31(.a2(a2[19:15]), .a3(a3[19:15]), .a4(a4[19:15]), .y(y1[19:15]));
	sbox_2 sb32(.a1(a1[19:15]), .a3(a3[19:15]), .a4(a4[19:15]), .y(y2[19:15]));
	sbox_3 sb33(.a1(a1[19:15]), .a2(a2[19:15]), .a4(a4[19:15]), .y(y3[19:15]));
	sbox_4 sb34(.a1(a1[19:15]), .a2(a2[19:15]), .a3(a3[19:15]), .y(y4[19:15]));

	sbox_1 sb41(.a2(a2[24:20]), .a3(a3[24:20]), .a4(a4[24:20]), .y(y1[24:20]));
	sbox_2 sb42(.a1(a1[24:20]), .a3(a3[24:20]), .a4(a4[24:20]), .y(y2[24:20]));
	sbox_3 sb43(.a1(a1[24:20]), .a2(a2[24:20]), .a4(a4[24:20]), .y(y3[24:20]));
	sbox_4 sb44(.a1(a1[24:20]), .a2(a2[24:20]), .a3(a3[24:20]), .y(y4[24:20]));

	sbox_1 sb51(.a2(a2[29:25]), .a3(a3[29:25]), .a4(a4[29:25]), .y(y1[29:25]));
	sbox_2 sb52(.a1(a1[29:25]), .a3(a3[29:25]), .a4(a4[29:25]), .y(y2[29:25]));
	sbox_3 sb53(.a1(a1[29:25]), .a2(a2[29:25]), .a4(a4[29:25]), .y(y3[29:25]));
	sbox_4 sb54(.a1(a1[29:25]), .a2(a2[29:25]), .a3(a3[29:25]), .y(y4[29:25]));

	sbox_1 sb61(.a2(a2[34:30]), .a3(a3[34:30]), .a4(a4[34:30]), .y(y1[34:30]));
	sbox_2 sb62(.a1(a1[34:30]), .a3(a3[34:30]), .a4(a4[34:30]), .y(y2[34:30]));
	sbox_3 sb63(.a1(a1[34:30]), .a2(a2[34:30]), .a4(a4[34:30]), .y(y3[34:30]));
	sbox_4 sb64(.a1(a1[34:30]), .a2(a2[34:30]), .a3(a3[34:30]), .y(y4[34:30]));

	sbox_1 sb71(.a2(a2[39:35]), .a3(a3[39:35]), .a4(a4[39:35]), .y(y1[39:35]));
	sbox_2 sb72(.a1(a1[39:35]), .a3(a3[39:35]), .a4(a4[39:35]), .y(y2[39:35]));
	sbox_3 sb73(.a1(a1[39:35]), .a2(a2[39:35]), .a4(a4[39:35]), .y(y3[39:35]));
	sbox_4 sb74(.a1(a1[39:35]), .a2(a2[39:35]), .a3(a3[39:35]), .y(y4[39:35]));

	sbox_1 sb81(.a2(a2[44:40]), .a3(a3[44:40]), .a4(a4[44:40]), .y(y1[44:40]));
	sbox_2 sb82(.a1(a1[44:40]), .a3(a3[44:40]), .a4(a4[44:40]), .y(y2[44:40]));
	sbox_3 sb83(.a1(a1[44:40]), .a2(a2[44:40]), .a4(a4[44:40]), .y(y3[44:40]));
	sbox_4 sb84(.a1(a1[44:40]), .a2(a2[44:40]), .a3(a3[44:40]), .y(y4[44:40]));

	sbox_1 sb91(.a2(a2[49:45]), .a3(a3[49:45]), .a4(a4[49:45]), .y(y1[49:45]));
	sbox_2 sb92(.a1(a1[49:45]), .a3(a3[49:45]), .a4(a4[49:45]), .y(y2[49:45]));
	sbox_3 sb93(.a1(a1[49:45]), .a2(a2[49:45]), .a4(a4[49:45]), .y(y3[49:45]));
	sbox_4 sb94(.a1(a1[49:45]), .a2(a2[49:45]), .a3(a3[49:45]), .y(y4[49:45]));

	sbox_1 sb101(.a2(a2[54:50]), .a3(a3[54:50]), .a4(a4[54:50]), .y(y1[54:50]));
	sbox_2 sb102(.a1(a1[54:50]), .a3(a3[54:50]), .a4(a4[54:50]), .y(y2[54:50]));
	sbox_3 sb103(.a1(a1[54:50]), .a2(a2[54:50]), .a4(a4[54:50]), .y(y3[54:50]));
	sbox_4 sb104(.a1(a1[54:50]), .a2(a2[54:50]), .a3(a3[54:50]), .y(y4[54:50]));

	sbox_1 sb111(.a2(a2[59:55]), .a3(a3[59:55]), .a4(a4[59:55]), .y(y1[59:55]));
	sbox_2 sb112(.a1(a1[59:55]), .a3(a3[59:55]), .a4(a4[59:55]), .y(y2[59:55]));
	sbox_3 sb113(.a1(a1[59:55]), .a2(a2[59:55]), .a4(a4[59:55]), .y(y3[59:55]));
	sbox_4 sb114(.a1(a1[59:55]), .a2(a2[59:55]), .a3(a3[59:55]), .y(y4[59:55]));

	sbox_1 sb121(.a2(a2[64:60]), .a3(a3[64:60]), .a4(a4[64:60]), .y(y1[64:60]));
	sbox_2 sb122(.a1(a1[64:60]), .a3(a3[64:60]), .a4(a4[64:60]), .y(y2[64:60]));
	sbox_3 sb123(.a1(a1[64:60]), .a2(a2[64:60]), .a4(a4[64:60]), .y(y3[64:60]));
	sbox_4 sb124(.a1(a1[64:60]), .a2(a2[64:60]), .a3(a3[64:60]), .y(y4[64:60]));

	sbox_1 sb131(.a2(a2[69:65]), .a3(a3[69:65]), .a4(a4[69:65]), .y(y1[69:65]));
	sbox_2 sb132(.a1(a1[69:65]), .a3(a3[69:65]), .a4(a4[69:65]), .y(y2[69:65]));
	sbox_3 sb133(.a1(a1[69:65]), .a2(a2[69:65]), .a4(a4[69:65]), .y(y3[69:65]));
	sbox_4 sb134(.a1(a1[69:65]), .a2(a2[69:65]), .a3(a3[69:65]), .y(y4[69:65]));

	sbox_1 sb141(.a2(a2[74:70]), .a3(a3[74:70]), .a4(a4[74:70]), .y(y1[74:70]));
	sbox_2 sb142(.a1(a1[74:70]), .a3(a3[74:70]), .a4(a4[74:70]), .y(y2[74:70]));
	sbox_3 sb143(.a1(a1[74:70]), .a2(a2[74:70]), .a4(a4[74:70]), .y(y3[74:70]));
	sbox_4 sb144(.a1(a1[74:70]), .a2(a2[74:70]), .a3(a3[74:70]), .y(y4[74:70]));

	sbox_1 sb151(.a2(a2[79:75]), .a3(a3[79:75]), .a4(a4[79:75]), .y(y1[79:75]));
	sbox_2 sb152(.a1(a1[79:75]), .a3(a3[79:75]), .a4(a4[79:75]), .y(y2[79:75]));
	sbox_3 sb153(.a1(a1[79:75]), .a2(a2[79:75]), .a4(a4[79:75]), .y(y3[79:75]));
	sbox_4 sb154(.a1(a1[79:75]), .a2(a2[79:75]), .a3(a3[79:75]), .y(y4[79:75]));

	sbox_1 sb161(.a2(a2[84:80]), .a3(a3[84:80]), .a4(a4[84:80]), .y(y1[84:80]));
	sbox_2 sb162(.a1(a1[84:80]), .a3(a3[84:80]), .a4(a4[84:80]), .y(y2[84:80]));
	sbox_3 sb163(.a1(a1[84:80]), .a2(a2[84:80]), .a4(a4[84:80]), .y(y3[84:80]));
	sbox_4 sb164(.a1(a1[84:80]), .a2(a2[84:80]), .a3(a3[84:80]), .y(y4[84:80]));

	sbox_1 sb171(.a2(a2[89:85]), .a3(a3[89:85]), .a4(a4[89:85]), .y(y1[89:85]));
	sbox_2 sb172(.a1(a1[89:85]), .a3(a3[89:85]), .a4(a4[89:85]), .y(y2[89:85]));
	sbox_3 sb173(.a1(a1[89:85]), .a2(a2[89:85]), .a4(a4[89:85]), .y(y3[89:85]));
	sbox_4 sb174(.a1(a1[89:85]), .a2(a2[89:85]), .a3(a3[89:85]), .y(y4[89:85]));

	sbox_1 sb181(.a2(a2[94:90]), .a3(a3[94:90]), .a4(a4[94:90]), .y(y1[94:90]));
	sbox_2 sb182(.a1(a1[94:90]), .a3(a3[94:90]), .a4(a4[94:90]), .y(y2[94:90]));
	sbox_3 sb183(.a1(a1[94:90]), .a2(a2[94:90]), .a4(a4[94:90]), .y(y3[94:90]));
	sbox_4 sb184(.a1(a1[94:90]), .a2(a2[94:90]), .a3(a3[94:90]), .y(y4[94:90]));

	sbox_1 sb191(.a2(a2[99:95]), .a3(a3[99:95]), .a4(a4[99:95]), .y(y1[99:95]));
	sbox_2 sb192(.a1(a1[99:95]), .a3(a3[99:95]), .a4(a4[99:95]), .y(y2[99:95]));
	sbox_3 sb193(.a1(a1[99:95]), .a2(a2[99:95]), .a4(a4[99:95]), .y(y3[99:95]));
	sbox_4 sb194(.a1(a1[99:95]), .a2(a2[99:95]), .a3(a3[99:95]), .y(y4[99:95]));

	sbox_1 sb201(.a2(a2[104:100]), .a3(a3[104:100]), .a4(a4[104:100]), .y(y1[104:100]));
	sbox_2 sb202(.a1(a1[104:100]), .a3(a3[104:100]), .a4(a4[104:100]), .y(y2[104:100]));
	sbox_3 sb203(.a1(a1[104:100]), .a2(a2[104:100]), .a4(a4[104:100]), .y(y3[104:100]));
	sbox_4 sb204(.a1(a1[104:100]), .a2(a2[104:100]), .a3(a3[104:100]), .y(y4[104:100]));

	sbox_1 sb211(.a2(a2[109:105]), .a3(a3[109:105]), .a4(a4[109:105]), .y(y1[109:105]));
	sbox_2 sb212(.a1(a1[109:105]), .a3(a3[109:105]), .a4(a4[109:105]), .y(y2[109:105]));
	sbox_3 sb213(.a1(a1[109:105]), .a2(a2[109:105]), .a4(a4[109:105]), .y(y3[109:105]));
	sbox_4 sb214(.a1(a1[109:105]), .a2(a2[109:105]), .a3(a3[109:105]), .y(y4[109:105]));

	sbox_1 sb221(.a2(a2[114:110]), .a3(a3[114:110]), .a4(a4[114:110]), .y(y1[114:110]));
	sbox_2 sb222(.a1(a1[114:110]), .a3(a3[114:110]), .a4(a4[114:110]), .y(y2[114:110]));
	sbox_3 sb223(.a1(a1[114:110]), .a2(a2[114:110]), .a4(a4[114:110]), .y(y3[114:110]));
	sbox_4 sb224(.a1(a1[114:110]), .a2(a2[114:110]), .a3(a3[114:110]), .y(y4[114:110]));

	sbox_1 sb231(.a2(a2[119:115]), .a3(a3[119:115]), .a4(a4[119:115]), .y(y1[119:115]));
	sbox_2 sb232(.a1(a1[119:115]), .a3(a3[119:115]), .a4(a4[119:115]), .y(y2[119:115]));
	sbox_3 sb233(.a1(a1[119:115]), .a2(a2[119:115]), .a4(a4[119:115]), .y(y3[119:115]));
	sbox_4 sb234(.a1(a1[119:115]), .a2(a2[119:115]), .a3(a3[119:115]), .y(y4[119:115]));

	sbox_1 sb241(.a2(a2[124:120]), .a3(a3[124:120]), .a4(a4[124:120]), .y(y1[124:120]));
	sbox_2 sb242(.a1(a1[124:120]), .a3(a3[124:120]), .a4(a4[124:120]), .y(y2[124:120]));
	sbox_3 sb243(.a1(a1[124:120]), .a2(a2[124:120]), .a4(a4[124:120]), .y(y3[124:120]));
	sbox_4 sb244(.a1(a1[124:120]), .a2(a2[124:120]), .a3(a3[124:120]), .y(y4[124:120]));

	sbox_1 sb251(.a2(a2[129:125]), .a3(a3[129:125]), .a4(a4[129:125]), .y(y1[129:125]));
	sbox_2 sb252(.a1(a1[129:125]), .a3(a3[129:125]), .a4(a4[129:125]), .y(y2[129:125]));
	sbox_3 sb253(.a1(a1[129:125]), .a2(a2[129:125]), .a4(a4[129:125]), .y(y3[129:125]));
	sbox_4 sb254(.a1(a1[129:125]), .a2(a2[129:125]), .a3(a3[129:125]), .y(y4[129:125]));

	sbox_1 sb261(.a2(a2[134:130]), .a3(a3[134:130]), .a4(a4[134:130]), .y(y1[134:130]));
	sbox_2 sb262(.a1(a1[134:130]), .a3(a3[134:130]), .a4(a4[134:130]), .y(y2[134:130]));
	sbox_3 sb263(.a1(a1[134:130]), .a2(a2[134:130]), .a4(a4[134:130]), .y(y3[134:130]));
	sbox_4 sb264(.a1(a1[134:130]), .a2(a2[134:130]), .a3(a3[134:130]), .y(y4[134:130]));

	sbox_1 sb271(.a2(a2[139:135]), .a3(a3[139:135]), .a4(a4[139:135]), .y(y1[139:135]));
	sbox_2 sb272(.a1(a1[139:135]), .a3(a3[139:135]), .a4(a4[139:135]), .y(y2[139:135]));
	sbox_3 sb273(.a1(a1[139:135]), .a2(a2[139:135]), .a4(a4[139:135]), .y(y3[139:135]));
	sbox_4 sb274(.a1(a1[139:135]), .a2(a2[139:135]), .a3(a3[139:135]), .y(y4[139:135]));

	sbox_1 sb281(.a2(a2[144:140]), .a3(a3[144:140]), .a4(a4[144:140]), .y(y1[144:140]));
	sbox_2 sb282(.a1(a1[144:140]), .a3(a3[144:140]), .a4(a4[144:140]), .y(y2[144:140]));
	sbox_3 sb283(.a1(a1[144:140]), .a2(a2[144:140]), .a4(a4[144:140]), .y(y3[144:140]));
	sbox_4 sb284(.a1(a1[144:140]), .a2(a2[144:140]), .a3(a3[144:140]), .y(y4[144:140]));

	sbox_1 sb291(.a2(a2[149:145]), .a3(a3[149:145]), .a4(a4[149:145]), .y(y1[149:145]));
	sbox_2 sb292(.a1(a1[149:145]), .a3(a3[149:145]), .a4(a4[149:145]), .y(y2[149:145]));
	sbox_3 sb293(.a1(a1[149:145]), .a2(a2[149:145]), .a4(a4[149:145]), .y(y3[149:145]));
	sbox_4 sb294(.a1(a1[149:145]), .a2(a2[149:145]), .a3(a3[149:145]), .y(y4[149:145]));

	sbox_1 sb301(.a2(a2[154:150]), .a3(a3[154:150]), .a4(a4[154:150]), .y(y1[154:150]));
	sbox_2 sb302(.a1(a1[154:150]), .a3(a3[154:150]), .a4(a4[154:150]), .y(y2[154:150]));
	sbox_3 sb303(.a1(a1[154:150]), .a2(a2[154:150]), .a4(a4[154:150]), .y(y3[154:150]));
	sbox_4 sb304(.a1(a1[154:150]), .a2(a2[154:150]), .a3(a3[154:150]), .y(y4[154:150]));

	sbox_1 sb311(.a2(a2[159:155]), .a3(a3[159:155]), .a4(a4[159:155]), .y(y1[159:155]));
	sbox_2 sb312(.a1(a1[159:155]), .a3(a3[159:155]), .a4(a4[159:155]), .y(y2[159:155]));
	sbox_3 sb313(.a1(a1[159:155]), .a2(a2[159:155]), .a4(a4[159:155]), .y(y3[159:155]));
	sbox_4 sb314(.a1(a1[159:155]), .a2(a2[159:155]), .a3(a3[159:155]), .y(y4[159:155]));

 endmodule 
